package reg_8bit_config;
	parameter R=8;
endpackage
