package Verilog_parameter;
parameter S = 8;
endpackage
