package v8_parameters;
parameter k=7;
parameter l=7;
parameter M=16;
endpackage 