package v11_filter_parameters;
	parameter	k = 8;
	parameter	l = 5;
	parameter	M = 16;
	parameter   N = 13; //k + l
endpackage