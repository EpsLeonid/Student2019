package q2par;
parameter Width = 8;
endpackage