package Zadanie2_parameter;
parameter R=8;
endpackage
