package v10_parameters;
parameter N_10=16;
parameter K_10=10;
parameter L_10=6;
parameter M_10=16;
endpackage

