package Task_2_5;
	parameter N = 8;
endpackage 