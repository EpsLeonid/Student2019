package Pollparametr;
parameter Const = 8;
endpackage