module proj_1

(
input wire operandA,
input wire operandB,
output wire out_mul
);



assign out_mul=operandA*operandB;

endmodule
