package v17_filter_parameters;	 
	parameter k_17	= 10;
	parameter l_17 = 5;
	parameter M_17	= 16;
	parameter N_17 = 15;
	parameter SizE = 20;
endpackage 