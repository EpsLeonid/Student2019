//������������ ������
package sun_parameter;
parameter sun=8;
endpackage
