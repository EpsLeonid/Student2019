package v15_filter_parameters;
	parameter	v15_k = 6;
	parameter	v15_l = 6;
	parameter	v15_M = 16;
	parameter 	v15_bufferSize = 13;
	parameter	v15_dataSize = 20;
endpackage
