package Zadanie_2_parameter;
parameter R = 8;
parameter outR = 16;
endpackage