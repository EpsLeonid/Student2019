package SysVerParam;
parameter P = 8;
endpackage