package v14_parameters;
parameter K_14=9;
parameter L_14=5;
parameter M_14=16;
endpackage
