package v15_filter_parameters;
	parameter	k = 6;
	parameter	l = 6;
	parameter	M = 16;
	parameter   T1 = 16;
	parameter   T2 = 5;
	parameter 	bufferSize = 12;
	parameter	dataSize = 20;
endpackage
