package ABC_parameter;
parameter WIDTH=8;
endpackage
