package v7_filter_parameters;

//Parameter declaration
parameter k = 10;
parameter l = 5;
parameter M = 5;

endpackage