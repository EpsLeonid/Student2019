package parameters;
	//файл с параметром, который определяет размер регистра
	parameter sizeOfReg = 8;
	
endpackage
