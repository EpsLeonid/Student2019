package V1_par;
parameter Const=8;
endpackage