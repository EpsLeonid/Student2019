module Task2(input A,B, output C);
	assign C=A*B;// ������ ������� � � � � �� ������������ � ����������� ������� �
endmodule