package v20_filter_param;

parameter k = 10;
parameter l = 6;
parameter M = 16;
parameter SIZE_ADC_DATA = 16;
parameter SIZE_REG = 16;
parameter SIZE_FILTER_DATA = 16;
endpackage