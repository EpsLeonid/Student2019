package v11_filter_parameters;
	parameter	k_11 = 8;
	parameter	l_11 = 5;
	parameter	M_11 = 16;
	parameter   N_11 = 13; //k + l
endpackage