package argum;
//����������� ����������� ��� 
parameter size=8;
parameter DATA_OUT_size=16;

endpackage 