package v3_parameters;

parameter k_3=11;
parameter l_3=5;
parameter m1_3=16;
parameter m2_3=1;
parameter SIZE = 20;
endpackage

