package v18_filter_parameters;	 
parameter k_19	= 7;
parameter l_19 = 7;
parameter M_19	= 16;
parameter N_19 = 15;
parameter MSize_19 = 20;
endpackage 