/*
	������� ������ ������������� � ��������,
	� ����� ��� �������������.
	������� �� ��������� ��������� �������� ������ ������������� �� ����

	��������� ������ D-��������.
*/
module AB
(
	// ���������� ������� ��������
	input A,
	input B,
	input clk,
	// ���������� �������� ��������
	output q
);

logic a,b; // �������� ��� �������� ������� �������� 
logic ab; // ������� �������� ������� A*B

// ������������ ������� ������
d_trigger dtrigA(.d(A),.clk(clk),.out(a)); 
d_trigger dtrigB(.d(B),.clk(clk),.out(b));


always_ff @(posedge clk) // �� ��������� ������ clk �������...
begin
	ab <= a * b;
end

assign q = ab; // ����������� ������

endmodule