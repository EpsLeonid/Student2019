package v14_parameters;
parameter N_14=13; //N_14=K_14+L_14
parameter K_14=9;
parameter L_14=5;
parameter M_14=16;
endpackage
