package v12_filter_parameters;
	parameter	m_12 = 16;
	parameter	k_12 = 5;
	parameter	l_12 = 5;
	parameter	size = 20;
	parameter	numSliceData = 10;
endpackage