package parameters;
	parameter	k = 5;
	parameter	l = 5;
	parameter	M = 16;
	parameter	numSliceData = 10;
	endpackage