package v19_parameters;
parameter L = 6;
parameter K = 13;
parameter M1 = 15;
parameter M2 = 1;
parameter memSize = 13;
endpackage
