//������������ ������
//������� ���������� �������

package v13_parameters;

	parameter l_13 = 5;
	parameter k_13 = 11;
	parameter m1 = 16;
	parameter m2 = 1;
	parameter SIZE = 20;
	
endpackage
