package Zadan_2_par;
parameter input_size = 8;
parameter outinput_size = 16;
endpackage