package v16_parameters;
parameter l_16 = 6;
parameter k_16 = 13;
parameter m1_16 = 16;
parameter m2_16 = 1;
parameter saveDataSize = 16;
endpackage