package testparametr;
parameter Width = 8;
endpackage