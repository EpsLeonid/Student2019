package v5_parameters;
parameter N_5=13; //N=K+L
parameter K_5=6;
parameter L_5=6;
parameter M_5=16;
endpackage
