package v1_parameters;
parameter N=13; //N=K+L
parameter K=8;
parameter L=5;
parameter M=16;
endpackage
