package v2_parameters;
parameter N_2=10; 
parameter K_2=5;
parameter L_2=5;
parameter M_2=16;
endpackage

