package v9_parameters;
parameter L = 6;
parameter K = 13;
parameter M1 = 15;
parameter M2 = 1;
parameter memSize1 = 13;
endpackage
