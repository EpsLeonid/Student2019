package module_2_parameter;
parameter par = 7;
endpackage
