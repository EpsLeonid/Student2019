//������������ ������
//������� ���������� �������


package v13_parameters;

	parameter l_13 = 5;
	parameter k_13 = 11;
	parameter N_13 = 16;
	parameter m1_13 = 16;
	parameter m2_13 = 1;
	parameter SIZE = 20;
	
	
endpackage
