package v19_parameters;
	parameter l_19 = 6;
	parameter k_19 = 13;
	parameter N_19 = 13;
	parameter m1_19 = 15;
	parameter m2_19 = 1;
	parameter SIZE19 = 20;
	
endpackage
