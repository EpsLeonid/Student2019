package v6_parameters;
parameter l_6 = 6;
parameter k_6 = 13;
parameter m1_6 = 16;
parameter m2_6 = 1;
parameter saveDataSize = 13;
endpackage