package v7_filter_parameters;

//Parameter declaration
parameter k_7 = 10;
parameter l_7 = 5;
parameter M_7 = 16;
parameter N_7 = 15;
parameter S_7 = 20;

endpackage