module multSignals(
	input signal_1,
	input signal_2,
	output mult
);
	assign mult=signal_1*signal_2;
endmodule
