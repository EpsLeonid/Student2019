package parameters;
	//���� � ����������, ������� ���������� ������ ��������
	parameter sizeOfReg = 8;
	
endpackage
