package v21_filter_parameters;
	parameter	v21_k = 5;
	parameter	v21_l = 5;
	parameter	v21_M = 15;
	parameter 	v21_array = 10; //k+l
	parameter	v21_Size = 20;
endpackage
