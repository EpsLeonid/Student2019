package v9_parameters;
	parameter l_9 = 6;
	parameter k_9 = 13;
	parameter N_9 = 13;
	parameter m1_9 = 15;
	parameter m2_9 = 1;
	parameter SIZE9 = 20;
	
endpackage