package parameters;
	// ����������� ������ ��� ������
	parameter	a_size = 8;
	parameter	b_size = 8;
	parameter	c_size = 8;
	parameter	data_size = a_size * 2;

endpackage 