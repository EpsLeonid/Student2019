package testparametr;
parameter Const = 8;
endpackage