package Task_25;
 parameter N=8;
endpackage