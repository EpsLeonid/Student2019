package v1_parameters;
parameter N_1=13; //N=K+L
parameter K_1=8;
parameter L_1=5;
parameter M_1=16;
endpackage
