//�������������� ������

package par_parameter;
parameter par = 7;

endpackage
