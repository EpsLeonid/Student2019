package module_2_1_parameter;
parameter katusha=8;
endpackage
