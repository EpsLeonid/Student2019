module Task_2_2(output C, input A, B);
	assign C = A & B;
endmodule 