package v12_filter_parameters;
	parameter	m = 16;
	parameter	k = 5;
	parameter	l = 5;
	parameter	size = 20;
	parameter	numSliceData = 10;
endpackage