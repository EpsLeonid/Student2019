package SystemVerilog1Param;
parameter P = 8;
endpackage