import module_2_parameter::par; // ����������� ����� � ����������

module module_2 
(
	// ������ ������� 2.2
	input wire a,
	input wire b,
	output wire c,
	
	// ������ ������� 2.3
	input clk,
	input d,
	output exit,
	
	//������ ������� 2.4
	input [par:0]A,
	input [par:0]B,
	input [par:0]C,
	output [par*2+1:0]out  
);
// ������� 2.2
assign c = b*a;
	
// ������� 2.3
always@(posedge clk) // �� ��������� ������ clk
begin
exit <=d;
end
	
// ������� 2.4
// �������� ��������� A1,B1,C1,C2	
reg [par:0]A1;
reg [par:0]B1;
reg [par:0]C1;
reg [par:0]C2;

// �������� �������������� �������� R ��� �������� ����������� ���������
reg [par*2+1:0]R;

// �������� �������� out_1 ��� �������� ������������� ����������
reg [par*2+1:0]out_1;

always@(posedge clk)
begin
	C1<=C; // ������ � � ������� C1, � ����� � �2 �� clk 
	C2<=C1;
	A1<=A; // ������ A � ������� A1 �� clk
	B1<=B; // ������ B � ������� B1 �� clk
	
	// ������ ����������� ��������� � R
	R<=A1*B1;
	// ������ ������������� ����������� ���������� � out_1
	out_1 <= R+C2;	
end	

assign out = out_1;

endmodule 